//////////////////////////////////////////////////////////////////////////////////
// Design: OR gate using MUX
// Engineer: kiran
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module or_mux(
    input  wire A,
    input  wire B,
    output wire Z
    );

    mux u1 (.A(B), .B(A), .Sel(A), .Z(Z));

endmodule
