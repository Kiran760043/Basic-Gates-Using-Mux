//////////////////////////////////////////////////////////////////////////////////
// Design: XOR gate using MUX 
// Engineer: kiran
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps


module xor_mux(
    input  wire A,
    input  wire B,
    output wire Z
    );

    mux u1 (.A(B), .B(~B), .Sel(A), .Z(Z));

endmodule
