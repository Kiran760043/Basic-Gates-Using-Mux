//////////////////////////////////////////////////////////////////////////////////
// Design: AND gate using MUX 
// Engineer: kiran
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module and_mux(
    input A,
    input B,
    output Z
    );
    
    mux u1 (.A(A), .B(B), .Sel(A), .Z(Z));
    
endmodule
